-- megafunction wizard: %ALTASMI_PARALLEL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTASMI_PARALLEL 

-- ============================================================
-- File Name: asmi.vhd
-- Megafunction Name(s):
-- 			ALTASMI_PARALLEL
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1.dp6 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altasmi_parallel CBX_AUTO_BLACKBOX="ALL" DATA_WIDTH="STANDARD" DEVICE_FAMILY="Cyclone IV E" EPCS_TYPE="EPCS64" PAGE_SIZE=1 PORT_BULK_ERASE="PORT_UNUSED" PORT_DIE_ERASE="PORT_UNUSED" PORT_EN4B_ADDR="PORT_UNUSED" PORT_FAST_READ="PORT_UNUSED" PORT_ILLEGAL_ERASE="PORT_UNUSED" PORT_ILLEGAL_WRITE="PORT_UNUSED" PORT_RDID_OUT="PORT_UNUSED" PORT_READ_ADDRESS="PORT_UNUSED" PORT_READ_DUMMYCLK="PORT_UNUSED" PORT_READ_RDID="PORT_UNUSED" PORT_READ_SID="PORT_UNUSED" PORT_READ_STATUS="PORT_UNUSED" PORT_SECTOR_ERASE="PORT_UNUSED" PORT_SECTOR_PROTECT="PORT_UNUSED" PORT_SHIFT_BYTES="PORT_UNUSED" PORT_WREN="PORT_UNUSED" PORT_WRITE="PORT_UNUSED" USE_ASMIBLOCK="OFF" USE_EAB="ON" WRITE_DUMMY_CLK=0 addr asmi_dataoe asmi_dataout asmi_dclk asmi_scein asmi_sdoin busy clkin data_valid dataout rden read reset INTENDED_DEVICE_FAMILY="Cyclone IV E" ALTERA_INTERNAL_OPTIONS=SUPPRESS_DA_RULE_INTERNAL=C106
--VERSION_BEGIN 13.0 cbx_a_gray2bin 2013:11:23:01:03:22:SJ cbx_a_graycounter 2013:11:23:01:03:22:SJ cbx_altasmi_parallel 2013:11:23:01:03:22:SJ cbx_altdpram 2013:11:23:01:03:22:SJ cbx_altsyncram 2013:11:23:01:03:22:SJ cbx_arriav 2013:11:23:01:03:22:SJ cbx_cyclone 2013:11:23:01:03:22:SJ cbx_cycloneii 2013:11:23:01:03:22:SJ cbx_fifo_common 2013:11:23:01:03:22:SJ cbx_lpm_add_sub 2013:11:23:01:03:22:SJ cbx_lpm_compare 2013:11:23:01:03:22:SJ cbx_lpm_counter 2013:11:23:01:03:23:SJ cbx_lpm_decode 2013:11:23:01:03:23:SJ cbx_lpm_mux 2013:11:23:01:03:23:SJ cbx_mgl 2013:11:23:01:10:57:SJ cbx_scfifo 2013:11:23:01:03:23:SJ cbx_stratix 2013:11:23:01:03:23:SJ cbx_stratixii 2013:11:23:01:03:23:SJ cbx_stratixiii 2013:11:23:01:03:23:SJ cbx_stratixv 2013:11:23:01:03:23:SJ cbx_util_mgl 2013:11:23:01:03:23:SJ  VERSION_END

 LIBRARY altera_mf;
 USE altera_mf.all;

--synthesis_resources = a_graycounter 3 lut 8 mux21 1 reg 66 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  asmi_altasmi_parallel_67k2 IS 
	 PORT 
	 ( 
		 addr	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 asmi_dataoe	:	OUT  STD_LOGIC;
		 asmi_dataout	:	IN  STD_LOGIC := '0';
		 asmi_dclk	:	OUT  STD_LOGIC;
		 asmi_scein	:	OUT  STD_LOGIC;
		 asmi_sdoin	:	OUT  STD_LOGIC;
		 busy	:	OUT  STD_LOGIC;
		 clkin	:	IN  STD_LOGIC;
		 data_valid	:	OUT  STD_LOGIC;
		 dataout	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 rden	:	IN  STD_LOGIC;
		 read	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0'
	 ); 
 END asmi_altasmi_parallel_67k2;

 ARCHITECTURE RTL OF asmi_altasmi_parallel_67k2 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "SUPPRESS_DA_RULE_INTERNAL=C106";

	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range133w138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_lg_w_q_range136w137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_clock	:	STD_LOGIC;
	 SIGNAL  wire_addbyte_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_end_operation85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addbyte_cntr_w_q_range133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range98w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_lg_w_q_range96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_in_operation25w26w27w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_end1_cyc_reg_in_wire28w29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_gen_cntr_w_q_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w296w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w91w293w294w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w91w298w299w300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w89w90w306w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w383w384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w293w294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w317w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w298w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w89w90w306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w93w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w91w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w91w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w91w298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w91w129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w91w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range87w92w109w110w111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range87w92w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_q_range88w89w90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range88w93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range88w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range87w92w109w110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range87w92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_lg_w_q_range88w89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_clk_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_w81w82w83w84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_stage_cntr_w_q_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_stage_cntr_w_q_range88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 add_msb_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_add_msb_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_addr_reg_d	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 addr_reg	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_addr_reg_ena	:	STD_LOGIC_VECTOR(23 DOWNTO 0);
	 SIGNAL  wire_addr_reg_w_q_range356w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 wire_asmi_opcode_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 asmi_opcode_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_asmi_opcode_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL  wire_asmi_opcode_reg_w_q_range143w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 busy_det_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 clr_read_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dffe2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 dvalid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_dvalid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_dvalid_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 dvalid_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end1_cyc_reg2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_hdlyreg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 end_rbyte_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_end_rbyte_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_end_rbyte_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 end_read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 ncs_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_ncs_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_ncs_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_ncs_reg_w_lg_q343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_read_data_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_data_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_data_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 wire_read_dout_reg_d	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 read_dout_reg	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_dout_reg_ena	:	STD_LOGIC_VECTOR(7 DOWNTO 0);
	 SIGNAL	 read_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 wire_read_reg_ena	:	STD_LOGIC;
	 SIGNAL	 shift_op_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage2_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage3_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 stage4_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	wire_mux211_dataout	:	STD_LOGIC;
	 SIGNAL  wire_w254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w197w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w190w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode154w155w156w238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode154w155w156w157w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w162w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode193w194w195w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode164w165w166w242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode164w165w166w167w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode186w187w188w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read322w323w324w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read370w437w438w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase39w379w380w381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode154w155w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode159w160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode169w174w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode169w174w175w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode169w170w244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode169w170w171w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode193w194w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode164w165w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode205w206w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode186w187w188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read322w323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read322w323w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read370w437w438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_sec_erase39w379w380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_4baddr146w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write177w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write48w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode148w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode148w149w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode179w248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode179w180w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode154w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode159w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode199w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode199w200w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode202w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode202w203w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode182w250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode182w183w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode210w262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode210w211w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode213w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode213w214w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode169w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode169w170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode164w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode205w206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode151w236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode151w152w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_load_opcode186w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage3_wire30w31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_start_poll308w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read322w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write57w104w105w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write57w58w371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read370w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_sec_erase39w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rden_wire375w376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie355w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_bulk_erase303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_nonvolatile289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_busy359w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_shift_opcode144w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage3_wire357w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_stage4_wire374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_start_poll308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write48w320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_addr_overdie453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_busy_wire1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_clkin_wire86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_fast_read321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_memadd388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_polling173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_rdid36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_volatile185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write_volatile192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_add_cycle68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_fast_read62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_ophdly24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_pgwr_data47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_end_read65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_rdid_wire7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_sid_wire6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_sec_protect_wire5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_st_busy_wire101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_pagewr_buf_not_empty_range53w54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode213w264w265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_load_opcode213w214w215w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w371w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_rden_wire375w376w377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy367w368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_busy359w360w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_stage4_wire406w407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode213w264w265w266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_load_opcode213w214w215w216w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_rden_wire375w376w377w378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_not_busy359w360w361w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w217w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w267w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w217w218w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w267w268w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w217w218w219w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w267w268w269w270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w217w218w219w220w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w267w268w269w270w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w217w218w219w220w221w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w267w268w269w270w271w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w217w218w219w220w221w222w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w223w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w273w274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w223w224w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w273w274w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w223w224w225w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w273w274w275w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w223w224w225w226w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w273w274w275w276w277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w223w224w225w226w227w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w273w274w275w276w277w278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w_lg_w223w224w225w226w227w228w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w229w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w229w230w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w126w127w128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w126w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read370w391w392w393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_do_read_sid122w123w124w125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read370w391w392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_sid122w123w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_read_stat401w402w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_do_write57w104w105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read370w405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read370w391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_sid122w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_read_stat401w402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write57w104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_do_write57w58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_data0out_wire409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_4baddr304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_sid122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_read_stat401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_sec_erase39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_wren305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_do_write57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_load_opcode281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rden_wire375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  addr_overdie :	STD_LOGIC;
	 SIGNAL  addr_overdie_pos :	STD_LOGIC;
	 SIGNAL  addr_reg_overdie :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  b4addr_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  berase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  busy_wire :	STD_LOGIC;
	 SIGNAL  clkin_wire :	STD_LOGIC;
	 SIGNAL  clr_addmsb_wire :	STD_LOGIC;
	 SIGNAL  clr_endrbyte_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire :	STD_LOGIC;
	 SIGNAL  clr_read_wire2 :	STD_LOGIC;
	 SIGNAL  clr_write_wire2 :	STD_LOGIC;
	 SIGNAL  data0out_wire :	STD_LOGIC;
	 SIGNAL  data_valid_wire :	STD_LOGIC;
	 SIGNAL  dataout_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  derase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  do_4baddr :	STD_LOGIC;
	 SIGNAL  do_bulk_erase :	STD_LOGIC;
	 SIGNAL  do_die_erase :	STD_LOGIC;
	 SIGNAL  do_fast_read :	STD_LOGIC;
	 SIGNAL  do_fread_epcq :	STD_LOGIC;
	 SIGNAL  do_freadwrv_polling :	STD_LOGIC;
	 SIGNAL  do_memadd :	STD_LOGIC;
	 SIGNAL  do_polling :	STD_LOGIC;
	 SIGNAL  do_read :	STD_LOGIC;
	 SIGNAL  do_read_nonvolatile :	STD_LOGIC;
	 SIGNAL  do_read_rdid :	STD_LOGIC;
	 SIGNAL  do_read_sid :	STD_LOGIC;
	 SIGNAL  do_read_stat :	STD_LOGIC;
	 SIGNAL  do_read_volatile :	STD_LOGIC;
	 SIGNAL  do_sec_erase :	STD_LOGIC;
	 SIGNAL  do_sec_prot :	STD_LOGIC;
	 SIGNAL  do_sprot_polling :	STD_LOGIC;
	 SIGNAL  do_wait_dummyclk :	STD_LOGIC;
	 SIGNAL  do_wren :	STD_LOGIC;
	 SIGNAL  do_write :	STD_LOGIC;
	 SIGNAL  do_write_polling :	STD_LOGIC;
	 SIGNAL  do_write_volatile :	STD_LOGIC;
	 SIGNAL  end1_cyc_gen_cntr_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_normal_in_wire :	STD_LOGIC;
	 SIGNAL  end1_cyc_reg_in_wire :	STD_LOGIC;
	 SIGNAL  end_add_cycle :	STD_LOGIC;
	 SIGNAL  end_add_cycle_mux_datab_wire :	STD_LOGIC;
	 SIGNAL  end_fast_read :	STD_LOGIC;
	 SIGNAL  end_one_cyc_pos :	STD_LOGIC;
	 SIGNAL  end_one_cycle :	STD_LOGIC;
	 SIGNAL  end_op_wire :	STD_LOGIC;
	 SIGNAL  end_operation :	STD_LOGIC;
	 SIGNAL  end_ophdly :	STD_LOGIC;
	 SIGNAL  end_pgwr_data :	STD_LOGIC;
	 SIGNAL  end_read :	STD_LOGIC;
	 SIGNAL  end_read_byte :	STD_LOGIC;
	 SIGNAL  fast_read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  freadwrv_sdoin :	STD_LOGIC;
	 SIGNAL  in_operation :	STD_LOGIC;
	 SIGNAL  load_opcode :	STD_LOGIC;
	 SIGNAL  memadd_sdoin :	STD_LOGIC;
	 SIGNAL  not_busy :	STD_LOGIC;
	 SIGNAL  oe_wire :	STD_LOGIC;
	 SIGNAL  pagewr_buf_not_empty :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  rden_wire :	STD_LOGIC;
	 SIGNAL  rdid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_data_reg_in_wire :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  read_rdid_wire :	STD_LOGIC;
	 SIGNAL  read_sid_wire :	STD_LOGIC;
	 SIGNAL  read_wire :	STD_LOGIC;
	 SIGNAL  rflagstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rnvdummyclk_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  rsid_sdoin :	STD_LOGIC;
	 SIGNAL  rstat_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  scein_wire :	STD_LOGIC;
	 SIGNAL  sdoin_wire :	STD_LOGIC;
	 SIGNAL  sec_protect_wire :	STD_LOGIC;
	 SIGNAL  secprot_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  secprot_sdoin :	STD_LOGIC;
	 SIGNAL  serase_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  shift_opcode :	STD_LOGIC;
	 SIGNAL  shift_opdata :	STD_LOGIC;
	 SIGNAL  shift_pgwr_data :	STD_LOGIC;
	 SIGNAL  st_busy_wire :	STD_LOGIC;
	 SIGNAL  stage2_wire :	STD_LOGIC;
	 SIGNAL  stage3_wire :	STD_LOGIC;
	 SIGNAL  stage4_wire :	STD_LOGIC;
	 SIGNAL  start_frpoll :	STD_LOGIC;
	 SIGNAL  start_poll :	STD_LOGIC;
	 SIGNAL  start_sppoll :	STD_LOGIC;
	 SIGNAL  start_wrpoll :	STD_LOGIC;
	 SIGNAL  to_sdoin_wire :	STD_LOGIC;
	 SIGNAL  wren_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wren_wire :	STD_LOGIC;
	 SIGNAL  write_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  write_prot_true :	STD_LOGIC;
	 SIGNAL  write_sdoin :	STD_LOGIC;
	 SIGNAL  wrvolatile_opcode :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_addr_range366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_range358w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_addr_reg_overdie_range354w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_b4addr_opcode_range145w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_berase_opcode_range153w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_dataout_wire_range408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_derase_opcode_range158w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_fast_read_opcode_range198w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_pagewr_buf_not_empty_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdid_opcode_range209w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rdummyclk_opcode_range191w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_read_opcode_range201w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rflagstat_opcode_range168w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rnvdummyclk_opcode_range181w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rsid_opcode_range212w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rstat_opcode_range172w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_secprot_opcode_range204w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_serase_opcode_range163w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wren_opcode_range150w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_write_opcode_range176w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_wrvolatile_opcode_range184w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 COMPONENT  a_graycounter
	 GENERIC 
	 (
		PVALUE	:	NATURAL := 0;
		WIDTH	:	NATURAL := 8;
		lpm_type	:	STRING := "a_graycounter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		q	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		qbin	:	OUT STD_LOGIC_VECTOR(width-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
 BEGIN

	wire_w254w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode193w194w195w196w(0) AND wire_w_rdummyclk_opcode_range253w(0);
	loop0 : FOR i IN 0 TO 6 GENERATE 
		wire_w197w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode193w194w195w196w(0) AND wire_w_rdummyclk_opcode_range191w(i);
	END GENERATE loop0;
	wire_w252w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode186w187w188w189w(0) AND wire_w_wrvolatile_opcode_range251w(0);
	loop1 : FOR i IN 0 TO 6 GENERATE 
		wire_w190w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode186w187w188w189w(0) AND wire_w_wrvolatile_opcode_range184w(i);
	END GENERATE loop1;
	wire_w440w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read370w437w438w439w(0) AND end_read_byte;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode154w155w156w238w(0) <= wire_w_lg_w_lg_w_lg_load_opcode154w155w156w(0) AND wire_w_berase_opcode_range237w(0);
	loop2 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode154w155w156w157w(i) <= wire_w_lg_w_lg_w_lg_load_opcode154w155w156w(0) AND wire_w_berase_opcode_range153w(i);
	END GENERATE loop2;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w240w(0) <= wire_w_lg_w_lg_w_lg_load_opcode159w160w161w(0) AND wire_w_derase_opcode_range239w(0);
	loop3 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w162w(i) <= wire_w_lg_w_lg_w_lg_load_opcode159w160w161w(0) AND wire_w_derase_opcode_range158w(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode193w194w195w196w(0) <= wire_w_lg_w_lg_w_lg_load_opcode193w194w195w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode164w165w166w242w(0) <= wire_w_lg_w_lg_w_lg_load_opcode164w165w166w(0) AND wire_w_serase_opcode_range241w(0);
	loop4 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode164w165w166w167w(i) <= wire_w_lg_w_lg_w_lg_load_opcode164w165w166w(0) AND wire_w_serase_opcode_range163w(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w260w(0) <= wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) AND wire_w_secprot_opcode_range259w(0);
	loop5 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(i) <= wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) AND wire_w_secprot_opcode_range204w(i);
	END GENERATE loop5;
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode186w187w188w189w(0) <= wire_w_lg_w_lg_w_lg_load_opcode186w187w188w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_read322w323w324w325w(0) <= wire_w_lg_w_lg_w_lg_do_read322w323w324w(0) AND end_one_cycle;
	wire_w_lg_w_lg_w_lg_w_lg_do_read370w437w438w439w(0) <= wire_w_lg_w_lg_w_lg_do_read370w437w438w(0) AND end_one_cyc_pos;
	wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase39w379w380w381w(0) <= wire_w_lg_w_lg_w_lg_do_sec_erase39w379w380w(0) AND end_operation;
	wire_w_lg_w_lg_w_lg_load_opcode154w155w156w(0) <= wire_w_lg_w_lg_load_opcode154w155w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_w_lg_load_opcode159w160w161w(0) <= wire_w_lg_w_lg_load_opcode159w160w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_w_lg_load_opcode169w174w246w(0) <= wire_w_lg_w_lg_load_opcode169w174w(0) AND wire_w_rstat_opcode_range245w(0);
	loop6 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode169w174w175w(i) <= wire_w_lg_w_lg_load_opcode169w174w(0) AND wire_w_rstat_opcode_range172w(i);
	END GENERATE loop6;
	wire_w_lg_w_lg_w_lg_load_opcode169w170w244w(0) <= wire_w_lg_w_lg_load_opcode169w170w(0) AND wire_w_rflagstat_opcode_range243w(0);
	loop7 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode169w170w171w(i) <= wire_w_lg_w_lg_load_opcode169w170w(0) AND wire_w_rflagstat_opcode_range168w(i);
	END GENERATE loop7;
	wire_w_lg_w_lg_w_lg_load_opcode193w194w195w(0) <= wire_w_lg_w_lg_load_opcode193w194w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_w_lg_load_opcode164w165w166w(0) <= wire_w_lg_w_lg_load_opcode164w165w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_w_lg_load_opcode205w206w207w(0) <= wire_w_lg_w_lg_load_opcode205w206w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_w_lg_load_opcode186w187w188w(0) <= wire_w_lg_w_lg_load_opcode186w187w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_w_lg_do_read322w323w324w(0) <= wire_w_lg_w_lg_do_read322w323w(0) AND wire_w_lg_w_lg_do_write48w320w(0);
	wire_w_lg_w_lg_w_lg_do_read322w323w382w(0) <= wire_w_lg_w_lg_do_read322w323w(0) AND clr_write_wire2;
	wire_w_lg_w_lg_w_lg_do_read370w437w438w(0) <= wire_w_lg_w_lg_do_read370w437w(0) AND wire_stage_cntr_w_lg_w_q_range87w92w(0);
	wire_w_lg_w_lg_w_lg_do_sec_erase39w379w380w(0) <= wire_w_lg_w_lg_do_sec_erase39w379w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_w_lg_do_4baddr146w147w(0) <= wire_w_lg_do_4baddr146w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_do_write177w178w(0) <= wire_w_lg_do_write177w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_do_write48w302w(0) <= wire_w_lg_do_write48w(0) AND end_pgwr_data;
	wire_w_lg_w_lg_load_opcode148w234w(0) <= wire_w_lg_load_opcode148w(0) AND wire_w_b4addr_opcode_range233w(0);
	loop8 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode148w149w(i) <= wire_w_lg_load_opcode148w(0) AND wire_w_b4addr_opcode_range145w(i);
	END GENERATE loop8;
	wire_w_lg_w_lg_load_opcode179w248w(0) <= wire_w_lg_load_opcode179w(0) AND wire_w_write_opcode_range247w(0);
	loop9 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode179w180w(i) <= wire_w_lg_load_opcode179w(0) AND wire_w_write_opcode_range176w(i);
	END GENERATE loop9;
	wire_w_lg_w_lg_load_opcode154w155w(0) <= wire_w_lg_load_opcode154w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_load_opcode159w160w(0) <= wire_w_lg_load_opcode159w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_load_opcode199w256w(0) <= wire_w_lg_load_opcode199w(0) AND wire_w_fast_read_opcode_range255w(0);
	loop10 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode199w200w(i) <= wire_w_lg_load_opcode199w(0) AND wire_w_fast_read_opcode_range198w(i);
	END GENERATE loop10;
	wire_w_lg_w_lg_load_opcode202w258w(0) <= wire_w_lg_load_opcode202w(0) AND wire_w_read_opcode_range257w(0);
	loop11 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode202w203w(i) <= wire_w_lg_load_opcode202w(0) AND wire_w_read_opcode_range201w(i);
	END GENERATE loop11;
	wire_w_lg_w_lg_load_opcode182w250w(0) <= wire_w_lg_load_opcode182w(0) AND wire_w_rnvdummyclk_opcode_range249w(0);
	loop12 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode182w183w(i) <= wire_w_lg_load_opcode182w(0) AND wire_w_rnvdummyclk_opcode_range181w(i);
	END GENERATE loop12;
	wire_w_lg_w_lg_load_opcode210w262w(0) <= wire_w_lg_load_opcode210w(0) AND wire_w_rdid_opcode_range261w(0);
	loop13 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode210w211w(i) <= wire_w_lg_load_opcode210w(0) AND wire_w_rdid_opcode_range209w(i);
	END GENERATE loop13;
	wire_w_lg_w_lg_load_opcode213w264w(0) <= wire_w_lg_load_opcode213w(0) AND wire_w_rsid_opcode_range263w(0);
	loop14 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode213w214w(i) <= wire_w_lg_load_opcode213w(0) AND wire_w_rsid_opcode_range212w(i);
	END GENERATE loop14;
	wire_w_lg_w_lg_load_opcode169w174w(0) <= wire_w_lg_load_opcode169w(0) AND wire_w_lg_do_polling173w(0);
	wire_w_lg_w_lg_load_opcode169w170w(0) <= wire_w_lg_load_opcode169w(0) AND do_polling;
	wire_w_lg_w_lg_load_opcode193w194w(0) <= wire_w_lg_load_opcode193w(0) AND wire_w_lg_do_write_volatile192w(0);
	wire_w_lg_w_lg_load_opcode164w165w(0) <= wire_w_lg_load_opcode164w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_load_opcode205w206w(0) <= wire_w_lg_load_opcode205w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_load_opcode151w236w(0) <= wire_w_lg_load_opcode151w(0) AND wire_w_wren_opcode_range235w(0);
	loop15 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_load_opcode151w152w(i) <= wire_w_lg_load_opcode151w(0) AND wire_w_wren_opcode_range150w(i);
	END GENERATE loop15;
	wire_w_lg_w_lg_load_opcode186w187w(0) <= wire_w_lg_load_opcode186w(0) AND wire_w_lg_do_read_volatile185w(0);
	wire_w_lg_w_lg_stage3_wire30w31w(0) <= wire_w_lg_stage3_wire30w(0) AND do_wait_dummyclk;
	wire_w_lg_w_lg_start_poll308w309w(0) <= wire_w_lg_start_poll308w(0) AND do_polling;
	wire_w_lg_w_lg_do_read322w323w(0) <= wire_w_lg_do_read322w(0) AND wire_w_lg_do_fast_read321w(0);
	wire_w_lg_w_lg_w_lg_w_lg_do_write57w104w105w106w(0) <= wire_w_lg_w_lg_w_lg_do_write57w104w105w(0) AND write_prot_true;
	wire_w_lg_w_lg_w_lg_do_write57w58w371w(0) <= wire_w_lg_w_lg_do_write57w58w(0) AND do_memadd;
	wire_w_lg_w_lg_do_read370w437w(0) <= wire_w_lg_do_read370w(0) AND wire_stage_cntr_w_q_range88w(0);
	wire_w_lg_w_lg_do_sec_erase39w379w(0) <= wire_w_lg_do_sec_erase39w(0) AND wire_w_lg_do_wren38w(0);
	wire_w_lg_w_lg_rden_wire375w376w(0) <= wire_w_lg_rden_wire375w(0) AND not_busy;
	wire_w_lg_addr_overdie365w(0) <= addr_overdie AND wire_w_addr_reg_overdie_range364w(0);
	loop16 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_addr_overdie355w(i) <= addr_overdie AND wire_w_addr_reg_overdie_range354w(i);
	END GENERATE loop16;
	wire_w_lg_do_4baddr146w(0) <= do_4baddr AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_do_bulk_erase303w(0) <= do_bulk_erase AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_do_read_nonvolatile289w(0) <= do_read_nonvolatile AND wire_addbyte_cntr_w_q_range133w(0);
	wire_w_lg_do_write177w(0) <= do_write AND wire_w_lg_do_read_stat37w(0);
	wire_w_lg_do_write55w(0) <= do_write AND wire_w_lg_w_pagewr_buf_not_empty_range53w54w(0);
	wire_w_lg_do_write48w(0) <= do_write AND shift_pgwr_data;
	wire_w_lg_load_opcode148w(0) <= load_opcode AND wire_w_lg_w_lg_do_4baddr146w147w(0);
	wire_w_lg_load_opcode179w(0) <= load_opcode AND wire_w_lg_w_lg_do_write177w178w(0);
	wire_w_lg_load_opcode154w(0) <= load_opcode AND do_bulk_erase;
	wire_w_lg_load_opcode159w(0) <= load_opcode AND do_die_erase;
	wire_w_lg_load_opcode199w(0) <= load_opcode AND do_fast_read;
	wire_w_lg_load_opcode202w(0) <= load_opcode AND do_read;
	wire_w_lg_load_opcode182w(0) <= load_opcode AND do_read_nonvolatile;
	wire_w_lg_load_opcode210w(0) <= load_opcode AND do_read_rdid;
	wire_w_lg_load_opcode213w(0) <= load_opcode AND do_read_sid;
	wire_w_lg_load_opcode169w(0) <= load_opcode AND do_read_stat;
	wire_w_lg_load_opcode193w(0) <= load_opcode AND do_read_volatile;
	wire_w_lg_load_opcode164w(0) <= load_opcode AND do_sec_erase;
	wire_w_lg_load_opcode205w(0) <= load_opcode AND do_sec_prot;
	wire_w_lg_load_opcode151w(0) <= load_opcode AND do_wren;
	wire_w_lg_load_opcode186w(0) <= load_opcode AND do_write_volatile;
	wire_w_lg_not_busy367w(0) <= not_busy AND wire_w_addr_range366w(0);
	loop17 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_not_busy359w(i) <= not_busy AND wire_w_addr_range358w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_shift_opcode144w(i) <= shift_opcode AND wire_asmi_opcode_reg_w_q_range143w(i);
	END GENERATE loop18;
	wire_w_lg_stage3_wire373w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w371w372w(0);
	wire_w_lg_stage3_wire404w(0) <= stage3_wire AND wire_w_lg_w_lg_w_lg_do_read_stat401w402w403w(0);
	wire_w_lg_stage3_wire40w(0) <= stage3_wire AND wire_w_lg_do_sec_erase39w(0);
	wire_w_lg_stage3_wire30w(0) <= stage3_wire AND do_fast_read;
	loop19 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_stage3_wire357w(i) <= stage3_wire AND wire_addr_reg_w_q_range356w(i);
	END GENERATE loop19;
	wire_w_lg_stage4_wire406w(0) <= stage4_wire AND wire_w_lg_w_lg_do_read370w405w(0);
	wire_w_lg_stage4_wire374w(0) <= stage4_wire AND addr_overdie;
	wire_w_lg_start_poll308w(0) <= start_poll AND do_read_stat;
	wire_w_lg_w_lg_do_write48w320w(0) <= NOT wire_w_lg_do_write48w(0);
	wire_w_lg_addr_overdie453w(0) <= NOT addr_overdie;
	wire_w_lg_busy_wire1w(0) <= NOT busy_wire;
	wire_w_lg_clkin_wire86w(0) <= NOT clkin_wire;
	wire_w_lg_do_fast_read321w(0) <= NOT do_fast_read;
	wire_w_lg_do_memadd388w(0) <= NOT do_memadd;
	wire_w_lg_do_polling173w(0) <= NOT do_polling;
	wire_w_lg_do_read322w(0) <= NOT do_read;
	wire_w_lg_do_read_rdid36w(0) <= NOT do_read_rdid;
	wire_w_lg_do_read_stat37w(0) <= NOT do_read_stat;
	wire_w_lg_do_read_volatile185w(0) <= NOT do_read_volatile;
	wire_w_lg_do_wren38w(0) <= NOT do_wren;
	wire_w_lg_do_write_volatile192w(0) <= NOT do_write_volatile;
	wire_w_lg_end_add_cycle68w(0) <= NOT end_add_cycle;
	wire_w_lg_end_fast_read62w(0) <= NOT end_fast_read;
	wire_w_lg_end_ophdly24w(0) <= NOT end_ophdly;
	wire_w_lg_end_pgwr_data47w(0) <= NOT end_pgwr_data;
	wire_w_lg_end_read65w(0) <= NOT end_read;
	wire_w_lg_rden_wire455w(0) <= NOT rden_wire;
	wire_w_lg_read_rdid_wire7w(0) <= NOT read_rdid_wire;
	wire_w_lg_read_sid_wire6w(0) <= NOT read_sid_wire;
	wire_w_lg_sec_protect_wire5w(0) <= NOT sec_protect_wire;
	wire_w_lg_st_busy_wire101w(0) <= NOT st_busy_wire;
	wire_w_lg_w_pagewr_buf_not_empty_range53w54w(0) <= NOT wire_w_pagewr_buf_not_empty_range53w(0);
	wire_w_lg_w_lg_w_lg_load_opcode213w264w265w(0) <= wire_w_lg_w_lg_load_opcode213w264w(0) OR wire_w_lg_w_lg_load_opcode210w262w(0);
	loop20 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_load_opcode213w214w215w(i) <= wire_w_lg_w_lg_load_opcode213w214w(i) OR wire_w_lg_w_lg_load_opcode210w211w(i);
	END GENERATE loop20;
	wire_w_lg_w_lg_w_lg_w_lg_do_write57w58w371w372w(0) <= wire_w_lg_w_lg_w_lg_do_write57w58w371w(0) OR wire_w_lg_do_read370w(0);
	wire_w_lg_w_lg_w_lg_rden_wire375w376w377w(0) <= wire_w_lg_w_lg_rden_wire375w376w(0) OR wire_w_lg_stage4_wire374w(0);
	wire_w_lg_w_lg_not_busy367w368w(0) <= wire_w_lg_not_busy367w(0) OR wire_w_lg_addr_overdie365w(0);
	loop21 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_not_busy359w360w(i) <= wire_w_lg_not_busy359w(i) OR wire_w_lg_stage3_wire357w(i);
	END GENERATE loop21;
	wire_w_lg_w_lg_stage4_wire406w407w(0) <= wire_w_lg_stage4_wire406w(0) OR wire_w_lg_stage3_wire404w(0);
	wire_w_lg_w_lg_w_lg_w_lg_load_opcode213w264w265w266w(0) <= wire_w_lg_w_lg_w_lg_load_opcode213w264w265w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w260w(0);
	loop22 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_load_opcode213w214w215w216w(i) <= wire_w_lg_w_lg_w_lg_load_opcode213w214w215w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode205w206w207w208w(i);
	END GENERATE loop22;
	wire_w_lg_w_lg_w_lg_w_lg_rden_wire375w376w377w378w(0) <= wire_w_lg_w_lg_w_lg_rden_wire375w376w377w(0) OR wire_w_lg_stage3_wire373w(0);
	loop23 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_lg_w_lg_not_busy359w360w361w(i) <= wire_w_lg_w_lg_not_busy359w360w(i) OR wire_w_lg_addr_overdie355w(i);
	END GENERATE loop23;
	wire_w267w(0) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode213w264w265w266w(0) OR wire_w_lg_w_lg_load_opcode202w258w(0);
	loop24 : FOR i IN 0 TO 6 GENERATE 
		wire_w217w(i) <= wire_w_lg_w_lg_w_lg_w_lg_load_opcode213w214w215w216w(i) OR wire_w_lg_w_lg_load_opcode202w203w(i);
	END GENERATE loop24;
	wire_w_lg_w267w268w(0) <= wire_w267w(0) OR wire_w_lg_w_lg_load_opcode199w256w(0);
	loop25 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w217w218w(i) <= wire_w217w(i) OR wire_w_lg_w_lg_load_opcode199w200w(i);
	END GENERATE loop25;
	wire_w_lg_w_lg_w267w268w269w(0) <= wire_w_lg_w267w268w(0) OR wire_w254w(0);
	loop26 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w217w218w219w(i) <= wire_w_lg_w217w218w(i) OR wire_w197w(i);
	END GENERATE loop26;
	wire_w_lg_w_lg_w_lg_w267w268w269w270w(0) <= wire_w_lg_w_lg_w267w268w269w(0) OR wire_w252w(0);
	loop27 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w217w218w219w220w(i) <= wire_w_lg_w_lg_w217w218w219w(i) OR wire_w190w(i);
	END GENERATE loop27;
	wire_w_lg_w_lg_w_lg_w_lg_w267w268w269w270w271w(0) <= wire_w_lg_w_lg_w_lg_w267w268w269w270w(0) OR wire_w_lg_w_lg_load_opcode182w250w(0);
	loop28 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w217w218w219w220w221w(i) <= wire_w_lg_w_lg_w_lg_w217w218w219w220w(i) OR wire_w_lg_w_lg_load_opcode182w183w(i);
	END GENERATE loop28;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w267w268w269w270w271w272w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w267w268w269w270w271w(0) OR wire_w_lg_w_lg_load_opcode179w248w(0);
	loop29 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w217w218w219w220w221w222w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w217w218w219w220w221w(i) OR wire_w_lg_w_lg_load_opcode179w180w(i);
	END GENERATE loop29;
	wire_w273w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w267w268w269w270w271w272w(0) OR wire_w_lg_w_lg_w_lg_load_opcode169w174w246w(0);
	loop30 : FOR i IN 0 TO 6 GENERATE 
		wire_w223w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w217w218w219w220w221w222w(i) OR wire_w_lg_w_lg_w_lg_load_opcode169w174w175w(i);
	END GENERATE loop30;
	wire_w_lg_w273w274w(0) <= wire_w273w(0) OR wire_w_lg_w_lg_w_lg_load_opcode169w170w244w(0);
	loop31 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w223w224w(i) <= wire_w223w(i) OR wire_w_lg_w_lg_w_lg_load_opcode169w170w171w(i);
	END GENERATE loop31;
	wire_w_lg_w_lg_w273w274w275w(0) <= wire_w_lg_w273w274w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode164w165w166w242w(0);
	loop32 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w223w224w225w(i) <= wire_w_lg_w223w224w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode164w165w166w167w(i);
	END GENERATE loop32;
	wire_w_lg_w_lg_w_lg_w273w274w275w276w(0) <= wire_w_lg_w_lg_w273w274w275w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w240w(0);
	loop33 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w223w224w225w226w(i) <= wire_w_lg_w_lg_w223w224w225w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode159w160w161w162w(i);
	END GENERATE loop33;
	wire_w_lg_w_lg_w_lg_w_lg_w273w274w275w276w277w(0) <= wire_w_lg_w_lg_w_lg_w273w274w275w276w(0) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode154w155w156w238w(0);
	loop34 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w223w224w225w226w227w(i) <= wire_w_lg_w_lg_w_lg_w223w224w225w226w(i) OR wire_w_lg_w_lg_w_lg_w_lg_load_opcode154w155w156w157w(i);
	END GENERATE loop34;
	wire_w_lg_w_lg_w_lg_w_lg_w_lg_w273w274w275w276w277w278w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w273w274w275w276w277w(0) OR wire_w_lg_w_lg_load_opcode151w236w(0);
	loop35 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w_lg_w_lg_w_lg_w_lg_w223w224w225w226w227w228w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w223w224w225w226w227w(i) OR wire_w_lg_w_lg_load_opcode151w152w(i);
	END GENERATE loop35;
	wire_w279w(0) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w273w274w275w276w277w278w(0) OR wire_w_lg_w_lg_load_opcode148w234w(0);
	loop36 : FOR i IN 0 TO 6 GENERATE 
		wire_w229w(i) <= wire_w_lg_w_lg_w_lg_w_lg_w_lg_w223w224w225w226w227w228w(i) OR wire_w_lg_w_lg_load_opcode148w149w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 6 GENERATE 
		wire_w_lg_w229w230w(i) <= wire_w229w(i) OR wire_w_lg_shift_opcode144w(i);
	END GENERATE loop37;
	wire_w_lg_w_lg_w126w127w128w(0) <= wire_w_lg_w126w127w(0) OR do_read_nonvolatile;
	wire_w_lg_w126w127w(0) <= wire_w126w(0) OR do_fast_read;
	wire_w126w(0) <= wire_w_lg_w_lg_w_lg_w_lg_do_read_sid122w123w124w125w(0) OR do_read;
	wire_w_lg_w_lg_w_lg_w_lg_do_read370w391w392w393w(0) <= wire_w_lg_w_lg_w_lg_do_read370w391w392w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_w_lg_do_read_sid122w123w124w125w(0) <= wire_w_lg_w_lg_w_lg_do_read_sid122w123w124w(0) OR do_read_rdid;
	wire_w_lg_w_lg_w_lg_do_read370w391w392w(0) <= wire_w_lg_w_lg_do_read370w391w(0) OR do_sec_erase;
	wire_w_lg_w_lg_w_lg_do_read_sid122w123w124w(0) <= wire_w_lg_w_lg_do_read_sid122w123w(0) OR do_die_erase;
	wire_w_lg_w_lg_w_lg_do_read_stat401w402w403w(0) <= wire_w_lg_w_lg_do_read_stat401w402w(0) OR do_read_nonvolatile;
	wire_w_lg_w_lg_w_lg_do_write57w104w105w(0) <= wire_w_lg_w_lg_do_write57w104w(0) OR do_die_erase;
	wire_w_lg_w_lg_do_read370w405w(0) <= wire_w_lg_do_read370w(0) OR do_read_sid;
	wire_w_lg_w_lg_do_read370w391w(0) <= wire_w_lg_do_read370w(0) OR do_write;
	wire_w_lg_w_lg_do_read_sid122w123w(0) <= wire_w_lg_do_read_sid122w(0) OR do_sec_erase;
	wire_w_lg_w_lg_do_read_stat401w402w(0) <= wire_w_lg_do_read_stat401w(0) OR do_read_volatile;
	wire_w_lg_w_lg_do_write57w104w(0) <= wire_w_lg_do_write57w(0) OR do_bulk_erase;
	wire_w_lg_w_lg_do_write57w58w(0) <= wire_w_lg_do_write57w(0) OR do_die_erase;
	wire_w_lg_data0out_wire409w(0) <= data0out_wire OR wire_w_dataout_wire_range408w(0);
	wire_w_lg_do_4baddr304w(0) <= do_4baddr OR wire_w_lg_do_bulk_erase303w(0);
	wire_w_lg_do_read370w(0) <= do_read OR do_fast_read;
	wire_w_lg_do_read_sid122w(0) <= do_read_sid OR do_write;
	wire_w_lg_do_read_stat401w(0) <= do_read_stat OR do_read_rdid;
	wire_w_lg_do_sec_erase39w(0) <= do_sec_erase OR do_die_erase;
	wire_w_lg_do_wren305w(0) <= do_wren OR wire_w_lg_do_4baddr304w(0);
	wire_w_lg_do_write57w(0) <= do_write OR do_sec_erase;
	wire_w_lg_load_opcode281w(0) <= load_opcode OR shift_opcode;
	wire_w_lg_rden_wire375w(0) <= rden_wire OR wren_wire;
	addr_overdie <= '0';
	addr_overdie_pos <= '0';
	addr_reg_overdie <= (OTHERS => '0');
	asmi_dataoe <= oe_wire;
	asmi_dclk <= clkin_wire;
	asmi_scein <= scein_wire;
	asmi_sdoin <= sdoin_wire;
	b4addr_opcode <= (OTHERS => '0');
	berase_opcode <= (OTHERS => '0');
	busy <= busy_wire;
	busy_wire <= (((((((((((((do_read_rdid OR do_read_sid) OR do_read) OR do_fast_read) OR do_write) OR do_sec_prot) OR do_read_stat) OR do_sec_erase) OR do_bulk_erase) OR do_die_erase) OR do_4baddr) OR do_read_volatile) OR do_fread_epcq) OR do_read_nonvolatile);
	clkin_wire <= clkin;
	clr_addmsb_wire <= ((wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w383w384w(0) OR wire_w_lg_w_lg_w_lg_do_read322w323w382w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_sec_erase39w379w380w381w(0));
	clr_endrbyte_wire <= ((((wire_w_lg_do_read370w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR clr_read_wire2);
	clr_read_wire <= clr_read_reg;
	clr_read_wire2 <= clr_read_reg2;
	clr_write_wire2 <= '0';
	data0out_wire <= asmi_dataout;
	data_valid <= data_valid_wire;
	data_valid_wire <= dvalid_reg2;
	dataout <= ( read_data_reg(7 DOWNTO 0));
	dataout_wire <= ( "0000");
	derase_opcode <= (OTHERS => '0');
	do_4baddr <= '0';
	do_bulk_erase <= '0';
	do_die_erase <= '0';
	do_fast_read <= '0';
	do_fread_epcq <= '0';
	do_freadwrv_polling <= '0';
	do_memadd <= '0';
	do_polling <= ((do_write_polling OR do_sprot_polling) OR do_freadwrv_polling);
	do_read <= (((wire_w_lg_read_rdid_wire7w(0) AND wire_w_lg_read_sid_wire6w(0)) AND wire_w_lg_sec_protect_wire5w(0)) AND read_wire);
	do_read_nonvolatile <= '0';
	do_read_rdid <= '0';
	do_read_sid <= '0';
	do_read_stat <= '0';
	do_read_volatile <= '0';
	do_sec_erase <= '0';
	do_sec_prot <= '0';
	do_sprot_polling <= '0';
	do_wait_dummyclk <= '0';
	do_wren <= '0';
	do_write <= '0';
	do_write_polling <= '0';
	do_write_volatile <= '0';
	end1_cyc_gen_cntr_wire <= (wire_gen_cntr_w_lg_w_q_range98w99w(0) AND (NOT wire_gen_cntr_q(0)));
	end1_cyc_normal_in_wire <= (((((((((wire_stage_cntr_w_lg_w_lg_w_q_range87w92w109w(0) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_q(1)) AND wire_gen_cntr_q(0)) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range87w92w109w110w111w(0)) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write57w104w105w106w(0)) OR wire_w_lg_do_write55w(0)) OR ((do_read_stat AND start_poll) AND wire_w_lg_st_busy_wire101w(0)));
	end1_cyc_reg_in_wire <= end1_cyc_normal_in_wire;
	end_add_cycle <= wire_mux211_dataout;
	end_add_cycle_mux_datab_wire <= (wire_addbyte_cntr_q(2) AND wire_addbyte_cntr_q(1));
	end_fast_read <= end_read_reg;
	end_one_cyc_pos <= end1_cyc_reg2;
	end_one_cycle <= end1_cyc_reg;
	end_op_wire <= (((((((((((wire_stage_cntr_w_lg_w_q_range88w93w(0) AND ((wire_w_lg_w_lg_w_lg_w_lg_do_read322w323w324w325w(0) OR (do_read AND end_read)) OR (do_fast_read AND end_fast_read))) OR (wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w317w318w(0) AND wire_w_lg_do_polling173w(0))) OR ((((((do_read_rdid AND end_one_cyc_pos) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) AND wire_addbyte_cntr_q(2)) AND wire_addbyte_cntr_q(1)) AND wire_addbyte_cntr_w_lg_w_q_range136w137w(0))) OR (wire_w_lg_w_lg_start_poll308w309w(0) AND wire_w_lg_st_busy_wire101w(0))) OR wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w89w90w306w307w(0)) OR wire_w_lg_w_lg_w_lg_w_lg_do_write57w104w105w106w(0)) OR wire_w_lg_w_lg_do_write48w302w(0)) OR wire_w_lg_do_write55w(0)) OR wire_stage_cntr_w301w(0)) OR wire_stage_cntr_w_lg_w296w297w(0)) OR (wire_stage_cntr_w_lg_w_lg_w_q_range88w91w291w(0) AND ((do_write_volatile OR do_read_volatile) OR wire_w_lg_do_read_nonvolatile289w(0))));
	end_operation <= end_op_reg;
	end_ophdly <= end_op_hdlyreg;
	end_pgwr_data <= '0';
	end_read <= end_read_reg;
	end_read_byte <= (end_rbyte_reg AND wire_w_lg_addr_overdie453w(0));
	fast_read_opcode <= (OTHERS => '0');
	freadwrv_sdoin <= '0';
	in_operation <= busy_wire;
	load_opcode <= ((((wire_stage_cntr_w_lg_w_q_range88w89w(0) AND wire_stage_cntr_w_lg_w_q_range87w92w(0)) AND (NOT wire_gen_cntr_q(2))) AND wire_gen_cntr_w_lg_w_q_range96w97w(0)) AND wire_gen_cntr_q(0));
	memadd_sdoin <= add_msb_reg;
	not_busy <= busy_det_reg;
	oe_wire <= '0';
	pagewr_buf_not_empty <= ( "1");
	rden_wire <= rden;
	rdid_opcode <= (OTHERS => '0');
	rdummyclk_opcode <= (OTHERS => '0');
	read_data_reg_in_wire <= ( read_dout_reg(7 DOWNTO 0));
	read_opcode <= "00000011";
	read_rdid_wire <= '0';
	read_sid_wire <= '0';
	read_wire <= read_reg;
	rflagstat_opcode <= (OTHERS => '0');
	rnvdummyclk_opcode <= (OTHERS => '0');
	rsid_opcode <= (OTHERS => '0');
	rsid_sdoin <= '0';
	rstat_opcode <= (OTHERS => '0');
	scein_wire <= wire_ncs_reg_w_lg_q343w(0);
	sdoin_wire <= to_sdoin_wire;
	sec_protect_wire <= '0';
	secprot_opcode <= (OTHERS => '0');
	secprot_sdoin <= '0';
	serase_opcode <= (OTHERS => '0');
	shift_opcode <= shift_op_reg;
	shift_opdata <= stage2_wire;
	shift_pgwr_data <= '0';
	st_busy_wire <= '0';
	stage2_wire <= stage2_reg;
	stage3_wire <= stage3_reg;
	stage4_wire <= stage4_reg;
	start_frpoll <= '0';
	start_poll <= ((start_wrpoll OR start_sppoll) OR start_frpoll);
	start_sppoll <= '0';
	start_wrpoll <= '0';
	to_sdoin_wire <= ((((((shift_opdata AND asmi_opcode_reg(7)) OR rsid_sdoin) OR memadd_sdoin) OR write_sdoin) OR secprot_sdoin) OR freadwrv_sdoin);
	wren_opcode <= (OTHERS => '0');
	wren_wire <= '1';
	write_opcode <= (OTHERS => '0');
	write_prot_true <= '0';
	write_sdoin <= '0';
	wrvolatile_opcode <= (OTHERS => '0');
	wire_w_addr_range366w(0) <= addr(0);
	wire_w_addr_range358w <= addr(23 DOWNTO 1);
	wire_w_addr_reg_overdie_range364w(0) <= addr_reg_overdie(0);
	wire_w_addr_reg_overdie_range354w <= addr_reg_overdie(23 DOWNTO 1);
	wire_w_b4addr_opcode_range233w(0) <= b4addr_opcode(0);
	wire_w_b4addr_opcode_range145w <= b4addr_opcode(7 DOWNTO 1);
	wire_w_berase_opcode_range237w(0) <= berase_opcode(0);
	wire_w_berase_opcode_range153w <= berase_opcode(7 DOWNTO 1);
	wire_w_dataout_wire_range408w(0) <= dataout_wire(1);
	wire_w_derase_opcode_range239w(0) <= derase_opcode(0);
	wire_w_derase_opcode_range158w <= derase_opcode(7 DOWNTO 1);
	wire_w_fast_read_opcode_range255w(0) <= fast_read_opcode(0);
	wire_w_fast_read_opcode_range198w <= fast_read_opcode(7 DOWNTO 1);
	wire_w_pagewr_buf_not_empty_range53w(0) <= pagewr_buf_not_empty(0);
	wire_w_rdid_opcode_range261w(0) <= rdid_opcode(0);
	wire_w_rdid_opcode_range209w <= rdid_opcode(7 DOWNTO 1);
	wire_w_rdummyclk_opcode_range253w(0) <= rdummyclk_opcode(0);
	wire_w_rdummyclk_opcode_range191w <= rdummyclk_opcode(7 DOWNTO 1);
	wire_w_read_opcode_range257w(0) <= read_opcode(0);
	wire_w_read_opcode_range201w <= read_opcode(7 DOWNTO 1);
	wire_w_rflagstat_opcode_range243w(0) <= rflagstat_opcode(0);
	wire_w_rflagstat_opcode_range168w <= rflagstat_opcode(7 DOWNTO 1);
	wire_w_rnvdummyclk_opcode_range249w(0) <= rnvdummyclk_opcode(0);
	wire_w_rnvdummyclk_opcode_range181w <= rnvdummyclk_opcode(7 DOWNTO 1);
	wire_w_rsid_opcode_range263w(0) <= rsid_opcode(0);
	wire_w_rsid_opcode_range212w <= rsid_opcode(7 DOWNTO 1);
	wire_w_rstat_opcode_range245w(0) <= rstat_opcode(0);
	wire_w_rstat_opcode_range172w <= rstat_opcode(7 DOWNTO 1);
	wire_w_secprot_opcode_range259w(0) <= secprot_opcode(0);
	wire_w_secprot_opcode_range204w <= secprot_opcode(7 DOWNTO 1);
	wire_w_serase_opcode_range241w(0) <= serase_opcode(0);
	wire_w_serase_opcode_range163w <= serase_opcode(7 DOWNTO 1);
	wire_w_wren_opcode_range235w(0) <= wren_opcode(0);
	wire_w_wren_opcode_range150w <= wren_opcode(7 DOWNTO 1);
	wire_w_write_opcode_range247w(0) <= write_opcode(0);
	wire_w_write_opcode_range176w <= write_opcode(7 DOWNTO 1);
	wire_w_wrvolatile_opcode_range251w(0) <= wrvolatile_opcode(0);
	wire_w_wrvolatile_opcode_range184w <= wrvolatile_opcode(7 DOWNTO 1);
	wire_addbyte_cntr_w_lg_w_q_range133w138w(0) <= wire_addbyte_cntr_w_q_range133w(0) AND wire_addbyte_cntr_w_lg_w_q_range136w137w(0);
	wire_addbyte_cntr_w_lg_w_q_range136w137w(0) <= NOT wire_addbyte_cntr_w_q_range136w(0);
	wire_addbyte_cntr_clk_en <= wire_stage_cntr_w132w(0);
	wire_stage_cntr_w132w(0) <= ((wire_stage_cntr_w_lg_w_lg_w_q_range88w91w129w(0) AND wire_w_lg_w_lg_w126w127w128w(0)) OR addr_overdie) OR end_operation;
	wire_addbyte_cntr_clock <= wire_w_lg_clkin_wire86w(0);
	wire_addbyte_cntr_sclr <= wire_w_lg_end_operation85w(0);
	wire_w_lg_end_operation85w(0) <= end_operation OR addr_overdie;
	wire_addbyte_cntr_w_q_range136w(0) <= wire_addbyte_cntr_q(0);
	wire_addbyte_cntr_w_q_range133w(0) <= wire_addbyte_cntr_q(1);
	addbyte_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_addbyte_cntr_clk_en,
		clock => wire_addbyte_cntr_clock,
		q => wire_addbyte_cntr_q,
		sclr => wire_addbyte_cntr_sclr
	  );
	wire_gen_cntr_w_lg_w_q_range98w99w(0) <= wire_gen_cntr_w_q_range98w(0) AND wire_gen_cntr_w_lg_w_q_range96w97w(0);
	wire_gen_cntr_w_lg_w_q_range96w97w(0) <= NOT wire_gen_cntr_w_q_range96w(0);
	wire_gen_cntr_clk_en <= wire_w_lg_w_lg_w_lg_in_operation25w26w27w(0);
	wire_w_lg_w_lg_w_lg_in_operation25w26w27w(0) <= ((in_operation AND wire_w_lg_end_ophdly24w(0)) OR do_wait_dummyclk) OR addr_overdie;
	wire_gen_cntr_sclr <= wire_w_lg_w_lg_end1_cyc_reg_in_wire28w29w(0);
	wire_w_lg_w_lg_end1_cyc_reg_in_wire28w29w(0) <= (end1_cyc_reg_in_wire OR addr_overdie) OR do_wait_dummyclk;
	wire_gen_cntr_w_q_range96w(0) <= wire_gen_cntr_q(1);
	wire_gen_cntr_w_q_range98w(0) <= wire_gen_cntr_q(2);
	gen_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 3
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_gen_cntr_clk_en,
		clock => clkin_wire,
		q => wire_gen_cntr_q,
		sclr => wire_gen_cntr_sclr
	  );
	wire_stage_cntr_w_lg_w296w297w(0) <= wire_stage_cntr_w296w(0) AND end_one_cycle;
	wire_stage_cntr_w296w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w91w293w294w295w(0) AND end_add_cycle;
	wire_stage_cntr_w301w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w91w298w299w300w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w91w293w294w295w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w293w294w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w91w298w299w300w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w298w299w(0) AND wire_w_lg_do_read_stat37w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range88w89w90w306w307w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w89w90w306w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w93w383w384w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range88w93w383w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w293w294w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range88w91w293w(0) AND wire_w_lg_do_wren38w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w317w318w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range88w91w317w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w91w298w299w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range88w91w298w(0) AND wire_w_lg_do_wren38w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range88w89w90w306w(0) <= wire_stage_cntr_w_lg_w_lg_w_q_range88w89w90w(0) AND wire_w_lg_do_wren305w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range88w93w383w(0) <= wire_stage_cntr_w_lg_w_q_range88w93w(0) AND end_add_cycle;
	wire_stage_cntr_w_lg_w_lg_w_q_range88w91w293w(0) <= wire_stage_cntr_w_lg_w_q_range88w91w(0) AND wire_w_lg_do_sec_erase39w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range88w91w317w(0) <= wire_stage_cntr_w_lg_w_q_range88w91w(0) AND do_read_stat;
	wire_stage_cntr_w_lg_w_lg_w_q_range88w91w298w(0) <= wire_stage_cntr_w_lg_w_q_range88w91w(0) AND do_sec_prot;
	wire_stage_cntr_w_lg_w_lg_w_q_range88w91w129w(0) <= wire_stage_cntr_w_lg_w_q_range88w91w(0) AND end_one_cyc_pos;
	wire_stage_cntr_w_lg_w_lg_w_q_range88w91w291w(0) <= wire_stage_cntr_w_lg_w_q_range88w91w(0) AND end_one_cycle;
	wire_stage_cntr_w_lg_w_lg_w_lg_w_lg_w_q_range87w92w109w110w111w(0) <= wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range87w92w109w110w(0) AND end1_cyc_gen_cntr_wire;
	wire_stage_cntr_w_lg_w_lg_w_q_range87w92w109w(0) <= wire_stage_cntr_w_lg_w_q_range87w92w(0) AND wire_stage_cntr_w_lg_w_q_range88w89w(0);
	wire_stage_cntr_w_lg_w_lg_w_q_range88w89w90w(0) <= wire_stage_cntr_w_lg_w_q_range88w89w(0) AND wire_stage_cntr_w_q_range87w(0);
	wire_stage_cntr_w_lg_w_q_range88w93w(0) <= wire_stage_cntr_w_q_range88w(0) AND wire_stage_cntr_w_lg_w_q_range87w92w(0);
	wire_stage_cntr_w_lg_w_q_range88w91w(0) <= wire_stage_cntr_w_q_range88w(0) AND wire_stage_cntr_w_q_range87w(0);
	wire_stage_cntr_w_lg_w_lg_w_lg_w_q_range87w92w109w110w(0) <= NOT wire_stage_cntr_w_lg_w_lg_w_q_range87w92w109w(0);
	wire_stage_cntr_w_lg_w_q_range87w92w(0) <= NOT wire_stage_cntr_w_q_range87w(0);
	wire_stage_cntr_w_lg_w_q_range88w89w(0) <= NOT wire_stage_cntr_w_q_range88w(0);
	wire_stage_cntr_clk_en <= wire_w_lg_w_lg_w_lg_w81w82w83w84w(0);
	wire_w_lg_w_lg_w_lg_w81w82w83w84w(0) <= (((((((((((((in_operation AND end_one_cycle) AND (NOT (stage3_wire AND wire_w_lg_end_add_cycle68w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_read65w(0)))) AND (NOT (stage4_wire AND wire_w_lg_end_fast_read62w(0)))) AND (NOT ((wire_w_lg_w_lg_do_write57w58w(0) OR do_bulk_erase) AND write_prot_true))) AND (NOT wire_w_lg_do_write55w(0))) AND (NOT (stage3_wire AND st_busy_wire))) AND (NOT (wire_w_lg_do_write48w(0) AND wire_w_lg_end_pgwr_data47w(0)))) AND (NOT (stage2_wire AND do_wren))) AND (NOT (((wire_w_lg_stage3_wire40w(0) AND wire_w_lg_do_wren38w(0)) AND wire_w_lg_do_read_stat37w(0)) AND wire_w_lg_do_read_rdid36w(0)))) AND (NOT (stage3_wire AND ((do_write_volatile OR do_read_volatile) OR do_read_nonvolatile)))) OR wire_w_lg_w_lg_stage3_wire30w31w(0)) OR addr_overdie) OR end_ophdly;
	wire_stage_cntr_sclr <= wire_w_lg_end_operation85w(0);
	wire_stage_cntr_w_q_range87w(0) <= wire_stage_cntr_q(0);
	wire_stage_cntr_w_q_range88w(0) <= wire_stage_cntr_q(1);
	stage_cntr :  a_graycounter
	  GENERIC MAP (
		WIDTH => 2
	  )
	  PORT MAP ( 
		aclr => reset,
		clk_en => wire_stage_cntr_clk_en,
		clock => clkin_wire,
		q => wire_stage_cntr_q,
		sclr => wire_stage_cntr_sclr
	  );
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN add_msb_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_add_msb_reg_ena = '1') THEN 
				IF (clr_addmsb_wire = '1') THEN add_msb_reg <= '0';
				ELSE add_msb_reg <= addr_reg(23);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_add_msb_reg_ena <= ((((wire_w_lg_w_lg_w_lg_w_lg_do_read370w391w392w393w(0) AND (NOT (wire_w_lg_w_lg_do_write57w58w(0) AND wire_w_lg_do_memadd388w(0)))) AND wire_stage_cntr_q(1)) AND wire_stage_cntr_q(0)) OR clr_addmsb_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(0) = '1') THEN addr_reg(0) <= wire_addr_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(1) = '1') THEN addr_reg(1) <= wire_addr_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(2) = '1') THEN addr_reg(2) <= wire_addr_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(3) = '1') THEN addr_reg(3) <= wire_addr_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(4) = '1') THEN addr_reg(4) <= wire_addr_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(5) = '1') THEN addr_reg(5) <= wire_addr_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(6) = '1') THEN addr_reg(6) <= wire_addr_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(7) = '1') THEN addr_reg(7) <= wire_addr_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(8) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(8) = '1') THEN addr_reg(8) <= wire_addr_reg_d(8);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(9) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(9) = '1') THEN addr_reg(9) <= wire_addr_reg_d(9);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(10) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(10) = '1') THEN addr_reg(10) <= wire_addr_reg_d(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(11) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(11) = '1') THEN addr_reg(11) <= wire_addr_reg_d(11);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(12) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(12) = '1') THEN addr_reg(12) <= wire_addr_reg_d(12);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(13) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(13) = '1') THEN addr_reg(13) <= wire_addr_reg_d(13);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(14) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(14) = '1') THEN addr_reg(14) <= wire_addr_reg_d(14);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(15) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(15) = '1') THEN addr_reg(15) <= wire_addr_reg_d(15);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(16) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(16) = '1') THEN addr_reg(16) <= wire_addr_reg_d(16);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(17) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(17) = '1') THEN addr_reg(17) <= wire_addr_reg_d(17);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(18) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(18) = '1') THEN addr_reg(18) <= wire_addr_reg_d(18);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(19) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(19) = '1') THEN addr_reg(19) <= wire_addr_reg_d(19);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(20) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(20) = '1') THEN addr_reg(20) <= wire_addr_reg_d(20);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(21) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(21) = '1') THEN addr_reg(21) <= wire_addr_reg_d(21);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(22) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(22) = '1') THEN addr_reg(22) <= wire_addr_reg_d(22);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN addr_reg(23) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_addr_reg_ena(23) = '1') THEN addr_reg(23) <= wire_addr_reg_d(23);
			END IF;
		END IF;
	END PROCESS;
	wire_addr_reg_d <= ( wire_w_lg_w_lg_w_lg_not_busy359w360w361w & wire_w_lg_w_lg_not_busy367w368w);
	loop38 : FOR i IN 0 TO 23 GENERATE
		wire_addr_reg_ena(i) <= wire_w_lg_w_lg_w_lg_w_lg_rden_wire375w376w377w378w(0);
	END GENERATE loop38;
	wire_addr_reg_w_q_range356w <= addr_reg(22 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(0) = '1') THEN asmi_opcode_reg(0) <= wire_asmi_opcode_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(1) = '1') THEN asmi_opcode_reg(1) <= wire_asmi_opcode_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(2) = '1') THEN asmi_opcode_reg(2) <= wire_asmi_opcode_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(3) = '1') THEN asmi_opcode_reg(3) <= wire_asmi_opcode_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(4) = '1') THEN asmi_opcode_reg(4) <= wire_asmi_opcode_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(5) = '1') THEN asmi_opcode_reg(5) <= wire_asmi_opcode_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(6) = '1') THEN asmi_opcode_reg(6) <= wire_asmi_opcode_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN asmi_opcode_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_asmi_opcode_reg_ena(7) = '1') THEN asmi_opcode_reg(7) <= wire_asmi_opcode_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_asmi_opcode_reg_d <= ( wire_w_lg_w229w230w & wire_w279w);
	loop39 : FOR i IN 0 TO 7 GENERATE
		wire_asmi_opcode_reg_ena(i) <= wire_w_lg_load_opcode281w(0);
	END GENERATE loop39;
	wire_asmi_opcode_reg_w_q_range143w <= asmi_opcode_reg(6 DOWNTO 0);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN busy_det_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN busy_det_reg <= wire_w_lg_busy_wire1w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN clr_read_reg <= ((do_read_sid OR do_sec_prot) OR end_operation);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN clr_read_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN clr_read_reg2 <= clr_read_reg;
		END IF;
	END PROCESS;
	dffe2 <= '0';
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_dvalid_reg_ena = '1') THEN 
				IF (wire_dvalid_reg_sclr = '1') THEN dvalid_reg <= '0';
				ELSE dvalid_reg <= (end_read_byte AND end_one_cyc_pos);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_dvalid_reg_ena <= wire_w_lg_do_read370w(0);
	wire_dvalid_reg_sclr <= (end_op_wire OR end_operation);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN dvalid_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN dvalid_reg2 <= dvalid_reg;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end1_cyc_reg <= end1_cyc_reg_in_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end1_cyc_reg2 <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end1_cyc_reg2 <= end_one_cycle;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_hdlyreg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_op_hdlyreg <= end_operation;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN end_op_reg <= end_op_wire;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_rbyte_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_end_rbyte_reg_ena = '1') THEN 
				IF (wire_end_rbyte_reg_sclr = '1') THEN end_rbyte_reg <= '0';
				ELSE end_rbyte_reg <= wire_w_lg_w_lg_w_lg_do_read370w437w438w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_end_rbyte_reg_ena <= ((wire_gen_cntr_w_lg_w_q_range98w99w(0) AND wire_gen_cntr_q(0)) OR clr_endrbyte_wire);
	wire_end_rbyte_reg_sclr <= (clr_endrbyte_wire OR addr_overdie);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN end_read_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN end_read_reg <= (((wire_w_lg_rden_wire455w(0) AND wire_w_lg_do_read370w(0)) AND data_valid_wire) AND end_read_byte);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN ncs_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_ncs_reg_ena = '1') THEN 
				IF (wire_ncs_reg_sclr = '1') THEN ncs_reg <= '0';
				ELSE ncs_reg <= '1';
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_ncs_reg_ena <= (((wire_stage_cntr_w_lg_w_lg_w_q_range88w89w90w(0) AND end_one_cyc_pos) OR addr_overdie_pos) OR end_operation);
	wire_ncs_reg_sclr <= (end_operation OR addr_overdie_pos);
	wire_ncs_reg_w_lg_q343w(0) <= NOT ncs_reg;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(0) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(0) = '1') THEN read_data_reg(0) <= wire_read_data_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(1) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(1) = '1') THEN read_data_reg(1) <= wire_read_data_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(2) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(2) = '1') THEN read_data_reg(2) <= wire_read_data_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(3) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(3) = '1') THEN read_data_reg(3) <= wire_read_data_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(4) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(4) = '1') THEN read_data_reg(4) <= wire_read_data_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(5) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(5) = '1') THEN read_data_reg(5) <= wire_read_data_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(6) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(6) = '1') THEN read_data_reg(6) <= wire_read_data_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_data_reg(7) <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_data_reg_ena(7) = '1') THEN read_data_reg(7) <= wire_read_data_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_data_reg_d <= ( read_data_reg_in_wire(7 DOWNTO 0));
	loop40 : FOR i IN 0 TO 7 GENERATE
		wire_read_data_reg_ena(i) <= wire_w440w(0);
	END GENERATE loop40;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(0) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(0) = '1') THEN read_dout_reg(0) <= wire_read_dout_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(1) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(1) = '1') THEN read_dout_reg(1) <= wire_read_dout_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(2) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(2) = '1') THEN read_dout_reg(2) <= wire_read_dout_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(3) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(3) = '1') THEN read_dout_reg(3) <= wire_read_dout_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(4) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(4) = '1') THEN read_dout_reg(4) <= wire_read_dout_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(5) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(5) = '1') THEN read_dout_reg(5) <= wire_read_dout_reg_d(5);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(6) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(6) = '1') THEN read_dout_reg(6) <= wire_read_dout_reg_d(6);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_dout_reg(7) <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN 
			IF (wire_read_dout_reg_ena(7) = '1') THEN read_dout_reg(7) <= wire_read_dout_reg_d(7);
			END IF;
		END IF;
	END PROCESS;
	wire_read_dout_reg_d <= ( read_dout_reg(6 DOWNTO 0) & wire_w_lg_data0out_wire409w);
	loop41 : FOR i IN 0 TO 7 GENERATE
		wire_read_dout_reg_ena(i) <= wire_w_lg_w_lg_stage4_wire406w407w(0);
	END GENERATE loop41;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN read_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN 
			IF (wire_read_reg_ena = '1') THEN 
				IF (clr_read_wire = '1') THEN read_reg <= '0';
				ELSE read_reg <= read;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_read_reg_ena <= ((wire_w_lg_busy_wire1w(0) AND rden_wire) OR clr_read_wire);
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN shift_op_reg <= '0';
		ELSIF (clkin_wire = '1' AND clkin_wire'event) THEN shift_op_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range88w89w90w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage2_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage2_reg <= wire_stage_cntr_w_lg_w_lg_w_q_range88w89w90w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage3_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage3_reg <= wire_stage_cntr_w_lg_w_q_range88w91w(0);
		END IF;
	END PROCESS;
	PROCESS (clkin_wire, reset)
	BEGIN
		IF (reset = '1') THEN stage4_reg <= '0';
		ELSIF (clkin_wire = '0' AND clkin_wire'event) THEN stage4_reg <= wire_stage_cntr_w_lg_w_q_range88w93w(0);
		END IF;
	END PROCESS;
	wire_mux211_dataout <= end_add_cycle_mux_datab_wire WHEN do_fast_read = '1'  ELSE wire_addbyte_cntr_w_lg_w_q_range133w138w(0);

 END RTL; --asmi_altasmi_parallel_67k2
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY asmi IS
	PORT
	(
		addr		: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
		asmi_dataout		: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
		clkin		: IN STD_LOGIC ;
		rden		: IN STD_LOGIC ;
		read		: IN STD_LOGIC ;
		reset		: IN STD_LOGIC ;
		asmi_dataoe		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		asmi_dclk		: OUT STD_LOGIC ;
		asmi_scein		: OUT STD_LOGIC ;
		asmi_sdoin		: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
		busy		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		dataout		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
END asmi;


ARCHITECTURE RTL OF asmi IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "ALTASMI_PARALLEL";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "data_width=STANDARD;epcs_type=EPCS64;intended_device_family=Cyclone IV E;lpm_hint=UNUSED;lpm_type=altasmi_parallel;page_size=1;port_bulk_erase=PORT_UNUSED;port_die_erase=PORT_UNUSED;port_en4b_addr=PORT_UNUSED;port_fast_read=PORT_UNUSED;port_illegal_erase=PORT_UNUSED;port_illegal_write=PORT_UNUSED;port_rdid_out=PORT_UNUSED;port_read_address=PORT_UNUSED;port_read_dummyclk=PORT_UNUSED;port_read_rdid=PORT_UNUSED;port_read_sid=PORT_UNUSED;port_read_status=PORT_UNUSED;port_sector_erase=PORT_UNUSED;port_sector_protect=PORT_UNUSED;port_shift_bytes=PORT_UNUSED;port_wren=PORT_UNUSED;port_write=PORT_UNUSED;use_asmiblock=OFF;use_eab=ON;write_dummy_clk=0;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC ;



	COMPONENT asmi_altasmi_parallel_67k2
	PORT (
			read	: IN STD_LOGIC ;
			clkin	: IN STD_LOGIC ;
			data_valid	: OUT STD_LOGIC ;
			rden	: IN STD_LOGIC ;
			asmi_sdoin	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			dataout	: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
			addr	: IN STD_LOGIC_VECTOR (23 DOWNTO 0);
			asmi_dataoe	: OUT STD_LOGIC_VECTOR (0 DOWNTO 0);
			asmi_dataout	: IN STD_LOGIC_VECTOR (0 DOWNTO 0);
			asmi_dclk	: OUT STD_LOGIC ;
			asmi_scein	: OUT STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			reset	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	data_valid    <= sub_wire0;
	asmi_sdoin    <= sub_wire1(0 DOWNTO 0);
	dataout    <= sub_wire2(7 DOWNTO 0);
	asmi_dataoe    <= sub_wire3(0 DOWNTO 0);
	asmi_dclk    <= sub_wire4;
	asmi_scein    <= sub_wire5;
	busy    <= sub_wire6;

	asmi_altasmi_parallel_67k2_component : asmi_altasmi_parallel_67k2
	PORT MAP (
		read => read,
		clkin => clkin,
		rden => rden,
		addr => addr,
		asmi_dataout => asmi_dataout,
		reset => reset,
		data_valid => sub_wire0,
		asmi_sdoin => sub_wire1,
		dataout => sub_wire2,
		asmi_dataoe => sub_wire3,
		asmi_dclk => sub_wire4,
		asmi_scein => sub_wire5,
		busy => sub_wire6
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: DATA_WIDTH STRING "STANDARD"
-- Retrieval info: CONSTANT: EPCS_TYPE STRING "EPCS64"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: LPM_HINT STRING "UNUSED"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altasmi_parallel"
-- Retrieval info: CONSTANT: PAGE_SIZE NUMERIC "1"
-- Retrieval info: CONSTANT: PORT_BULK_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_DIE_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_EN4B_ADDR STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_FAST_READ STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_ILLEGAL_WRITE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_RDID_OUT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_ADDRESS STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_DUMMYCLK STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_RDID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_SID STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_READ_STATUS STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SECTOR_ERASE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SECTOR_PROTECT STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SHIFT_BYTES STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WREN STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_WRITE STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: USE_ASMIBLOCK STRING "OFF"
-- Retrieval info: CONSTANT: USE_EAB STRING "ON"
-- Retrieval info: CONSTANT: WRITE_DUMMY_CLK NUMERIC "0"
-- Retrieval info: USED_PORT: addr 0 0 24 0 INPUT NODEFVAL "addr[23..0]"
-- Retrieval info: CONNECT: @addr 0 0 24 0 addr 0 0 24 0
-- Retrieval info: USED_PORT: asmi_dataoe 0 0 1 0 OUTPUT NODEFVAL "asmi_dataoe[0..0]"
-- Retrieval info: CONNECT: asmi_dataoe 0 0 1 0 @asmi_dataoe 0 0 1 0
-- Retrieval info: USED_PORT: asmi_dataout 0 0 1 0 INPUT NODEFVAL "asmi_dataout[0..0]"
-- Retrieval info: CONNECT: @asmi_dataout 0 0 1 0 asmi_dataout 0 0 1 0
-- Retrieval info: USED_PORT: asmi_dclk 0 0 0 0 OUTPUT NODEFVAL "asmi_dclk"
-- Retrieval info: CONNECT: asmi_dclk 0 0 0 0 @asmi_dclk 0 0 0 0
-- Retrieval info: USED_PORT: asmi_scein 0 0 0 0 OUTPUT NODEFVAL "asmi_scein"
-- Retrieval info: CONNECT: asmi_scein 0 0 0 0 @asmi_scein 0 0 0 0
-- Retrieval info: USED_PORT: asmi_sdoin 0 0 1 0 OUTPUT NODEFVAL "asmi_sdoin[0..0]"
-- Retrieval info: CONNECT: asmi_sdoin 0 0 1 0 @asmi_sdoin 0 0 1 0
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: USED_PORT: clkin 0 0 0 0 INPUT NODEFVAL "clkin"
-- Retrieval info: CONNECT: @clkin 0 0 0 0 clkin 0 0 0 0
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: USED_PORT: dataout 0 0 8 0 OUTPUT NODEFVAL "dataout[7..0]"
-- Retrieval info: CONNECT: dataout 0 0 8 0 @dataout 0 0 8 0
-- Retrieval info: USED_PORT: rden 0 0 0 0 INPUT NODEFVAL "rden"
-- Retrieval info: CONNECT: @rden 0 0 0 0 rden 0 0 0 0
-- Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
-- Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
-- Retrieval info: USED_PORT: reset 0 0 0 0 INPUT NODEFVAL "reset"
-- Retrieval info: CONNECT: @reset 0 0 0 0 reset 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmi.vhd TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmi.qip TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmi.bsf FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmi_inst.vhd TRUE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmi.inc FALSE TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL asmi.cmp TRUE TRUE
